module to