module checker

import kdl.ast

fn kdl_parse_time(s string) {
}
