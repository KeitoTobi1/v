module kdl

pub type Any = Null
	| Time
	| DateTime
	| Date
	| i8
	| u8
	| i16
	| u16
	| int
	| u32
	| i64
	| u64
	| f32
	| f64
	| string

pub struct Date {
}

pub struct Time {
}

pub struct DateTime {
}
