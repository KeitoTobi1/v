// Copyright (c) 2024 Keito Tobichi All rights reserved.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.
module scanner

pub const next_line = rune(0x0085)
pub const form_feed = rune(0x000C)
pub const line_sep = rune(0x2028)
pub const paragraph_sep = rune(0x2029)
