module to

