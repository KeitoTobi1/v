// Copyright (c) 2024 Keito Tobichi All rights reserved.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.
module kdl

pub struct Null {
}

// decoding KDL Document.
pub fn decode(kdl_txt string) {
}

fn decode_struct() {
}

// parsing KDL query.
pub fn parse_query(query string) {
}

pub struct Uuid {
pub:
	uuid string
}

pub struct Uuidv6 {
pub:
	uuid_v6 string
}
